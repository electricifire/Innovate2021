-- mem_GN.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity mem_GN is
	port (
		Vbcont_int : out std_logic_vector(11 downto 0);        -- Vbcont_int.wire
		Clock      : in  std_logic                     := '0'; --      Clock.clk
		aclr       : in  std_logic                     := '0'; --           .reset_n
		Ibcont_int : out std_logic_vector(11 downto 0);        -- Ibcont_int.wire
		clk60KPLL  : in  std_logic                     := '0'; --  clk60KPLL.wire
		Iccont_int : out std_logic_vector(11 downto 0);        -- Iccont_int.wire
		Iacont_int : out std_logic_vector(11 downto 0);        -- Iacont_int.wire
		Vacont_int : out std_logic_vector(11 downto 0);        -- Vacont_int.wire
		Vccont_int : out std_logic_vector(11 downto 0)         -- Vccont_int.wire
	);
end entity mem_GN;

architecture rtl of mem_GN is
	component alt_dspbuilder_clock_GNF343OQUJ is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNF343OQUJ;

	component alt_dspbuilder_port_GN4K6H3QBP is
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN4K6H3QBP;

	component alt_dspbuilder_comparator_GN is
		generic (
			Operator  : string  := "Altaeb";
			lpm_width : natural := 8
		);
		port (
			clock  : in  std_logic                              := 'X';             -- clk
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			datab  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic;                                                 -- wire
			sclr   : in  std_logic                              := 'X'              -- clk
		);
	end component alt_dspbuilder_comparator_GN;

	component mem_GN_mem_Conversion_Ioxcont_Int1 is
		port (
			Ibcont     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			Iacont     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			Iacont_int : out std_logic_vector(12 downto 0);                    -- wire
			Ibcont_int : out std_logic_vector(12 downto 0);                    -- wire
			Clock      : in  std_logic                     := 'X';             -- clk
			aclr       : in  std_logic                     := 'X';             -- reset
			Iccont     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			Iccont_int : out std_logic_vector(12 downto 0)                     -- wire
		);
	end component mem_GN_mem_Conversion_Ioxcont_Int1;

	component alt_dspbuilder_rom_GNK7TUJIQA is
		generic (
			ClockPhase                : string   := "1";
			numwords                  : positive := 3;
			use_ena                   : natural  := 0;
			XFILE                     : string   := "input.hex";
			family                    : string   := "STRATIX";
			runtime_mod_instance_name : string   := "AAAA";
			register_outputs          : natural  := 1;
			data_width                : positive := 8;
			supportROM                : natural  := 1;
			ram_block_type            : string   := "AUTO";
			enable_runtime_mod        : natural  := 0;
			initialization            : string   := "From HEX file"
		);
		port (
			clock : in  std_logic                     := 'X';             -- clk
			aclr  : in  std_logic                     := 'X';             -- reset
			addr  : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- wire
			ena   : in  std_logic                     := 'X';             -- wire
			q     : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_rom_GNK7TUJIQA;

	component alt_dspbuilder_rom_GNLZO3EIT7 is
		generic (
			ClockPhase                : string   := "1";
			numwords                  : positive := 3;
			use_ena                   : natural  := 0;
			XFILE                     : string   := "input.hex";
			family                    : string   := "STRATIX";
			runtime_mod_instance_name : string   := "AAAA";
			register_outputs          : natural  := 1;
			data_width                : positive := 8;
			supportROM                : natural  := 1;
			ram_block_type            : string   := "AUTO";
			enable_runtime_mod        : natural  := 0;
			initialization            : string   := "From HEX file"
		);
		port (
			clock : in  std_logic                     := 'X';             -- clk
			aclr  : in  std_logic                     := 'X';             -- reset
			addr  : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- wire
			ena   : in  std_logic                     := 'X';             -- wire
			q     : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_rom_GNLZO3EIT7;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_constant_GN6XEGEZIQ is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(9 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN6XEGEZIQ;

	component mem_GN_mem_Conversion_Ioxcont_Int is
		port (
			vbcont     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			Vacont_int : out std_logic_vector(12 downto 0);                    -- wire
			Vbcont_int : out std_logic_vector(12 downto 0);                    -- wire
			Clock      : in  std_logic                     := 'X';             -- clk
			aclr       : in  std_logic                     := 'X';             -- reset
			vccont     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			vacont     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			Vccont_int : out std_logic_vector(12 downto 0)                     -- wire
		);
	end component mem_GN_mem_Conversion_Ioxcont_Int;

	component alt_dspbuilder_counter_GNWUDKEMTG is
		generic (
			svalue       : string  := "0";
			use_cnt_ena  : string  := "false";
			use_cout     : string  := "false";
			modulus      : integer := 256;
			use_sclr     : string  := "false";
			ndirection   : natural := 1;
			use_usr_aclr : string  := "false";
			width        : natural := 8;
			use_ena      : string  := "false";
			use_sset     : string  := "false";
			use_aload    : string  := "false";
			avalue       : string  := "0";
			use_aset     : string  := "false";
			use_sload    : string  := "false";
			use_cin      : string  := "false"
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			aload     : in  std_logic                          := 'X';             -- wire
			aset      : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cnt_ena   : in  std_logic                          := 'X';             -- wire
			cout      : out std_logic;                                             -- wire
			data      : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			direction : in  std_logic                          := 'X';             -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			q         : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr      : in  std_logic                          := 'X';             -- wire
			sload     : in  std_logic                          := 'X';             -- wire
			sset      : in  std_logic                          := 'X';             -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_counter_GNWUDKEMTG;

	component alt_dspbuilder_rom_GNOXA7UMVD is
		generic (
			ClockPhase                : string   := "1";
			numwords                  : positive := 3;
			use_ena                   : natural  := 0;
			XFILE                     : string   := "input.hex";
			family                    : string   := "STRATIX";
			runtime_mod_instance_name : string   := "AAAA";
			register_outputs          : natural  := 1;
			data_width                : positive := 8;
			supportROM                : natural  := 1;
			ram_block_type            : string   := "AUTO";
			enable_runtime_mod        : natural  := 0;
			initialization            : string   := "From HEX file"
		);
		port (
			clock : in  std_logic                     := 'X';             -- clk
			aclr  : in  std_logic                     := 'X';             -- reset
			addr  : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- wire
			ena   : in  std_logic                     := 'X';             -- wire
			q     : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_rom_GNOXA7UMVD;

	component alt_dspbuilder_cast_GN5D52DF5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- wire
			output : out std_logic_vector(10 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5D52DF5S;

	component alt_dspbuilder_cast_GNUDBRONP6 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(12 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNUDBRONP6;

	signal comparator1_result_wire                       : std_logic;                     -- Comparator1:result -> Counter1:sclr
	signal counter1_q_wire                               : std_logic_vector(9 downto 0);  -- Counter1:q -> [Sin1:addr, Sin2:addr, Sin:addr, cast79:input]
	signal sin_q_wire                                    : std_logic_vector(13 downto 0); -- Sin:q -> [mem_Conversion_Ioxcont_Int1_0:Iacont, mem_Conversion_Ioxcont_Int_0:vacont]
	signal sin1_q_wire                                   : std_logic_vector(13 downto 0); -- Sin1:q -> [mem_Conversion_Ioxcont_Int1_0:Ibcont, mem_Conversion_Ioxcont_Int_0:vbcont]
	signal sin2_q_wire                                   : std_logic_vector(13 downto 0); -- Sin2:q -> [mem_Conversion_Ioxcont_Int1_0:Iccont, mem_Conversion_Ioxcont_Int_0:vccont]
	signal clk60kpll_0_output_wire                       : std_logic;                     -- clk60KPLL_0:output -> [Counter1:ena, Sin1:ena, Sin2:ena, Sin:ena]
	signal constant2_output_wire                         : std_logic_vector(9 downto 0);  -- Constant2:output -> cast78:input
	signal cast78_output_wire                            : std_logic_vector(10 downto 0); -- cast78:output -> Comparator1:datab
	signal cast79_output_wire                            : std_logic_vector(10 downto 0); -- cast79:output -> Comparator1:dataa
	signal mem_conversion_ioxcont_int1_0_iacont_int_wire : std_logic_vector(12 downto 0); -- mem_Conversion_Ioxcont_Int1_0:Iacont_int -> cast80:input
	signal cast80_output_wire                            : std_logic_vector(11 downto 0); -- cast80:output -> Iacont_int_0:input
	signal mem_conversion_ioxcont_int1_0_ibcont_int_wire : std_logic_vector(12 downto 0); -- mem_Conversion_Ioxcont_Int1_0:Ibcont_int -> cast81:input
	signal cast81_output_wire                            : std_logic_vector(11 downto 0); -- cast81:output -> Ibcont_int_0:input
	signal mem_conversion_ioxcont_int1_0_iccont_int_wire : std_logic_vector(12 downto 0); -- mem_Conversion_Ioxcont_Int1_0:Iccont_int -> cast82:input
	signal cast82_output_wire                            : std_logic_vector(11 downto 0); -- cast82:output -> Iccont_int_0:input
	signal mem_conversion_ioxcont_int_0_vacont_int_wire  : std_logic_vector(12 downto 0); -- mem_Conversion_Ioxcont_Int_0:Vacont_int -> cast83:input
	signal cast83_output_wire                            : std_logic_vector(11 downto 0); -- cast83:output -> Vacont_int_0:input
	signal mem_conversion_ioxcont_int_0_vbcont_int_wire  : std_logic_vector(12 downto 0); -- mem_Conversion_Ioxcont_Int_0:Vbcont_int -> cast84:input
	signal cast84_output_wire                            : std_logic_vector(11 downto 0); -- cast84:output -> Vbcont_int_0:input
	signal mem_conversion_ioxcont_int_0_vccont_int_wire  : std_logic_vector(12 downto 0); -- mem_Conversion_Ioxcont_Int_0:Vccont_int -> cast85:input
	signal cast85_output_wire                            : std_logic_vector(11 downto 0); -- cast85:output -> Vccont_int_0:input
	signal clock_0_clock_output_clk                      : std_logic;                     -- Clock_0:clock_out -> [Comparator1:clock, Counter1:clock, Sin1:clock, Sin2:clock, Sin:clock, mem_Conversion_Ioxcont_Int1_0:Clock, mem_Conversion_Ioxcont_Int_0:Clock]
	signal clock_0_clock_output_reset                    : std_logic;                     -- Clock_0:aclr_out -> [Comparator1:sclr, Counter1:aclr, Sin1:aclr, Sin2:aclr, Sin:aclr, mem_Conversion_Ioxcont_Int1_0:aclr, mem_Conversion_Ioxcont_Int_0:aclr]

begin

	clock_0 : component alt_dspbuilder_clock_GNF343OQUJ
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr_n    => aclr                        --             .reset_n
		);

	iccont_int_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => cast82_output_wire, --  input.wire
			output => Iccont_int          -- output.wire
		);

	ibcont_int_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => cast81_output_wire, --  input.wire
			output => Ibcont_int          -- output.wire
		);

	comparator1 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altaeb",
			lpm_width => 11
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => cast79_output_wire,         --      dataa.wire
			datab  => cast78_output_wire,         --      datab.wire
			result => comparator1_result_wire     --     result.wire
		);

	iacont_int_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => cast80_output_wire, --  input.wire
			output => Iacont_int          -- output.wire
		);

	mem_conversion_ioxcont_int1_0 : component mem_GN_mem_Conversion_Ioxcont_Int1
		port map (
			Ibcont     => sin1_q_wire,                                   --     Ibcont.wire
			Iacont     => sin_q_wire,                                    --     Iacont.wire
			Iacont_int => mem_conversion_ioxcont_int1_0_iacont_int_wire, -- Iacont_int.wire
			Ibcont_int => mem_conversion_ioxcont_int1_0_ibcont_int_wire, -- Ibcont_int.wire
			Clock      => clock_0_clock_output_clk,                      --      Clock.clk
			aclr       => clock_0_clock_output_reset,                    --           .reset
			Iccont     => sin2_q_wire,                                   --     Iccont.wire
			Iccont_int => mem_conversion_ioxcont_int1_0_iccont_int_wire  -- Iccont_int.wire
		);

	sin2 : component alt_dspbuilder_rom_GNK7TUJIQA
		generic map (
			ClockPhase                => "1",
			numwords                  => 1000,
			use_ena                   => 1,
			XFILE                     => "input.hex",
			family                    => "Cyclone V",
			runtime_mod_instance_name => "AAAA",
			register_outputs          => 0,
			data_width                => 14,
			supportROM                => 1,
			ram_block_type            => "AUTO",
			enable_runtime_mod        => 0,
			initialization            => "From MATLAB array"
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			addr  => counter1_q_wire,            --       addr.wire
			ena   => clk60kpll_0_output_wire,    --        ena.wire
			q     => sin2_q_wire                 --          q.wire
		);

	sin1 : component alt_dspbuilder_rom_GNLZO3EIT7
		generic map (
			ClockPhase                => "1",
			numwords                  => 1000,
			use_ena                   => 1,
			XFILE                     => "input.hex",
			family                    => "Cyclone V",
			runtime_mod_instance_name => "AAAA",
			register_outputs          => 0,
			data_width                => 14,
			supportROM                => 1,
			ram_block_type            => "AUTO",
			enable_runtime_mod        => 0,
			initialization            => "From MATLAB array"
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			addr  => counter1_q_wire,            --       addr.wire
			ena   => clk60kpll_0_output_wire,    --        ena.wire
			q     => sin1_q_wire                 --          q.wire
		);

	clk60kpll_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => clk60KPLL,               --  input.wire
			output => clk60kpll_0_output_wire  -- output.wire
		);

	vccont_int_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => cast85_output_wire, --  input.wire
			output => Vccont_int          -- output.wire
		);

	vbcont_int_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => cast84_output_wire, --  input.wire
			output => Vbcont_int          -- output.wire
		);

	constant2 : component alt_dspbuilder_constant_GN6XEGEZIQ
		generic map (
			BitPattern => "1111101000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 10
		)
		port map (
			output => constant2_output_wire  -- output.wire
		);

	vacont_int_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => cast83_output_wire, --  input.wire
			output => Vacont_int          -- output.wire
		);

	mem_conversion_ioxcont_int_0 : component mem_GN_mem_Conversion_Ioxcont_Int
		port map (
			vbcont     => sin1_q_wire,                                  --     vbcont.wire
			Vacont_int => mem_conversion_ioxcont_int_0_vacont_int_wire, -- Vacont_int.wire
			Vbcont_int => mem_conversion_ioxcont_int_0_vbcont_int_wire, -- Vbcont_int.wire
			Clock      => clock_0_clock_output_clk,                     --      Clock.clk
			aclr       => clock_0_clock_output_reset,                   --           .reset
			vccont     => sin2_q_wire,                                  --     vccont.wire
			vacont     => sin_q_wire,                                   --     vacont.wire
			Vccont_int => mem_conversion_ioxcont_int_0_vccont_int_wire  -- Vccont_int.wire
		);

	counter1 : component alt_dspbuilder_counter_GNWUDKEMTG
		generic map (
			svalue       => "300",
			use_cnt_ena  => "false",
			use_cout     => "false",
			modulus      => 1000,
			use_sclr     => "true",
			ndirection   => 1,
			use_usr_aclr => "false",
			width        => 10,
			use_ena      => "true",
			use_sset     => "false",
			use_aload    => "false",
			avalue       => "0",
			use_aset     => "false",
			use_sload    => "false",
			use_cin      => "false"
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			ena   => clk60kpll_0_output_wire,    --        ena.wire
			sclr  => comparator1_result_wire,    --       sclr.wire
			q     => counter1_q_wire,            --          q.wire
			cout  => open                        --       cout.wire
		);

	sin : component alt_dspbuilder_rom_GNOXA7UMVD
		generic map (
			ClockPhase                => "1",
			numwords                  => 1000,
			use_ena                   => 1,
			XFILE                     => "input.hex",
			family                    => "Cyclone V",
			runtime_mod_instance_name => "AAAA",
			register_outputs          => 0,
			data_width                => 14,
			supportROM                => 1,
			ram_block_type            => "AUTO",
			enable_runtime_mod        => 0,
			initialization            => "From MATLAB array"
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			addr  => counter1_q_wire,            --       addr.wire
			ena   => clk60kpll_0_output_wire,    --        ena.wire
			q     => sin_q_wire                  --          q.wire
		);

	cast78 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant2_output_wire, --  input.wire
			output => cast78_output_wire     -- output.wire
		);

	cast79 : component alt_dspbuilder_cast_GN5D52DF5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter1_q_wire,    --  input.wire
			output => cast79_output_wire  -- output.wire
		);

	cast80 : component alt_dspbuilder_cast_GNUDBRONP6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => mem_conversion_ioxcont_int1_0_iacont_int_wire, --  input.wire
			output => cast80_output_wire                             -- output.wire
		);

	cast81 : component alt_dspbuilder_cast_GNUDBRONP6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => mem_conversion_ioxcont_int1_0_ibcont_int_wire, --  input.wire
			output => cast81_output_wire                             -- output.wire
		);

	cast82 : component alt_dspbuilder_cast_GNUDBRONP6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => mem_conversion_ioxcont_int1_0_iccont_int_wire, --  input.wire
			output => cast82_output_wire                             -- output.wire
		);

	cast83 : component alt_dspbuilder_cast_GNUDBRONP6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => mem_conversion_ioxcont_int_0_vacont_int_wire, --  input.wire
			output => cast83_output_wire                            -- output.wire
		);

	cast84 : component alt_dspbuilder_cast_GNUDBRONP6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => mem_conversion_ioxcont_int_0_vbcont_int_wire, --  input.wire
			output => cast84_output_wire                            -- output.wire
		);

	cast85 : component alt_dspbuilder_cast_GNUDBRONP6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => mem_conversion_ioxcont_int_0_vccont_int_wire, --  input.wire
			output => cast85_output_wire                            -- output.wire
		);

end architecture rtl; -- of mem_GN
