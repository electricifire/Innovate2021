-- mem_GN_mem_Conversion_Ioxcont_Int.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity mem_GN_mem_Conversion_Ioxcont_Int is
	port (
		vbcont     : in  std_logic_vector(13 downto 0) := (others => '0'); --     vbcont.wire
		Vacont_int : out std_logic_vector(12 downto 0);                    -- Vacont_int.wire
		Vbcont_int : out std_logic_vector(12 downto 0);                    -- Vbcont_int.wire
		Clock      : in  std_logic                     := '0';             --      Clock.clk
		aclr       : in  std_logic                     := '0';             --           .reset
		vccont     : in  std_logic_vector(13 downto 0) := (others => '0'); --     vccont.wire
		vacont     : in  std_logic_vector(13 downto 0) := (others => '0'); --     vacont.wire
		Vccont_int : out std_logic_vector(12 downto 0)                     -- Vccont_int.wire
	);
end entity mem_GN_mem_Conversion_Ioxcont_Int;

architecture rtl of mem_GN_mem_Conversion_Ioxcont_Int is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_multiplexer_GNBGHTTLA2 is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(12 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(12 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(12 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNBGHTTLA2;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_comparator_GN is
		generic (
			Operator  : string  := "Altaeb";
			lpm_width : natural := 8
		);
		port (
			clock  : in  std_logic                              := 'X';             -- clk
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			datab  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic;                                                 -- wire
			sclr   : in  std_logic                              := 'X'              -- clk
		);
	end component alt_dspbuilder_comparator_GN;

	component alt_dspbuilder_cast_GNUYRTQ4QH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNUYRTQ4QH;

	component alt_dspbuilder_pipelined_adder_GN4HTUTWRG is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GN4HTUTWRG;

	component alt_dspbuilder_constant_GN2SAWFEVT is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(12 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN2SAWFEVT;

	component alt_dspbuilder_constant_GNC5QUYE2B is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(12 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNC5QUYE2B;

	component alt_dspbuilder_cast_GN32Z4PX3B is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(30 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(30 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN32Z4PX3B;

	component alt_dspbuilder_constant_GNCOTI3HOF is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(10 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNCOTI3HOF;

	component alt_dspbuilder_constant_GNGPCXCFCV is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(12 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNGPCXCFCV;

	component alt_dspbuilder_cast_GNA5AA6QPF is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(12 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(12 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNA5AA6QPF;

	component alt_dspbuilder_port_GNBOOX3JQY is
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBOOX3JQY;

	component alt_dspbuilder_port_GNKZFR37ZH is
		port (
			input  : in  std_logic_vector(12 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(12 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNKZFR37ZH;

	component alt_dspbuilder_round_GNJN4GDIEL is
		generic (
			OUT_WIDTH_g     : natural := 6;
			IN_WIDTH_g      : natural := 8;
			PIPELINE_g      : natural := 0;
			ROUNDING_TYPE_g : string  := "TRUNCATE_LOW";
			SIGNED_g        : natural := 1
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- wire
			datain    : in  std_logic_vector(30 downto 0) := (others => 'X'); -- wire
			dataout   : out std_logic_vector(12 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_round_GNJN4GDIEL;

	component alt_dspbuilder_cast_GNVPCKFRV6 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNVPCKFRV6;

	component alt_dspbuilder_cast_GNL533AQU2 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(30 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNL533AQU2;

	component alt_dspbuilder_cast_GNSQKJ6AEZ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(30 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNSQKJ6AEZ;

	component alt_dspbuilder_cast_GND23XTBOL is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(30 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GND23XTBOL;

	component alt_dspbuilder_cast_GNRYH7CSLF is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(30 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNRYH7CSLF;

	component alt_dspbuilder_cast_GND5VHVYOD is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(30 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GND5VHVYOD;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	component alt_dspbuilder_cast_GNWF56JAW3 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(12 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNWF56JAW3;

	signal multiplexeruser_aclrgnd_output_wire       : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire             : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal pipelined_adder9user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder9user_aclrGND:output -> Pipelined_Adder9:user_aclr
	signal pipelined_adder9enavcc_output_wire        : std_logic;                     -- Pipelined_Adder9enaVCC:output -> Pipelined_Adder9:ena
	signal pipelined_adder4user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder4user_aclrGND:output -> Pipelined_Adder4:user_aclr
	signal pipelined_adder4enavcc_output_wire        : std_logic;                     -- Pipelined_Adder4enaVCC:output -> Pipelined_Adder4:ena
	signal pipelined_adder3user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder3user_aclrGND:output -> Pipelined_Adder3:user_aclr
	signal pipelined_adder3enavcc_output_wire        : std_logic;                     -- Pipelined_Adder3enaVCC:output -> Pipelined_Adder3:ena
	signal pipelined_adder2user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder2user_aclrGND:output -> Pipelined_Adder2:user_aclr
	signal pipelined_adder2enavcc_output_wire        : std_logic;                     -- Pipelined_Adder2enaVCC:output -> Pipelined_Adder2:ena
	signal pipelined_adder1user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder1user_aclrGND:output -> Pipelined_Adder1:user_aclr
	signal pipelined_adder1enavcc_output_wire        : std_logic;                     -- Pipelined_Adder1enaVCC:output -> Pipelined_Adder1:ena
	signal pipelined_adder8user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder8user_aclrGND:output -> Pipelined_Adder8:user_aclr
	signal pipelined_adder8enavcc_output_wire        : std_logic;                     -- Pipelined_Adder8enaVCC:output -> Pipelined_Adder8:ena
	signal pipelined_adder7user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder7user_aclrGND:output -> Pipelined_Adder7:user_aclr
	signal pipelined_adder7enavcc_output_wire        : std_logic;                     -- Pipelined_Adder7enaVCC:output -> Pipelined_Adder7:ena
	signal pipelined_adder6user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder6user_aclrGND:output -> Pipelined_Adder6:user_aclr
	signal pipelined_adder6enavcc_output_wire        : std_logic;                     -- Pipelined_Adder6enaVCC:output -> Pipelined_Adder6:ena
	signal pipelined_adder5user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder5user_aclrGND:output -> Pipelined_Adder5:user_aclr
	signal pipelined_adder5enavcc_output_wire        : std_logic;                     -- Pipelined_Adder5enaVCC:output -> Pipelined_Adder5:ena
	signal round1user_aclrgnd_output_wire            : std_logic;                     -- Round1user_aclrGND:output -> Round1:user_aclr
	signal round1enavcc_output_wire                  : std_logic;                     -- Round1enaVCC:output -> Round1:ena
	signal round1resetgnd_output_wire                : std_logic;                     -- Round1resetGND:output -> Round1:reset
	signal multiplexer3user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer3user_aclrGND:output -> Multiplexer3:user_aclr
	signal multiplexer3enavcc_output_wire            : std_logic;                     -- Multiplexer3enaVCC:output -> Multiplexer3:ena
	signal round2user_aclrgnd_output_wire            : std_logic;                     -- Round2user_aclrGND:output -> Round2:user_aclr
	signal round2enavcc_output_wire                  : std_logic;                     -- Round2enaVCC:output -> Round2:ena
	signal round2resetgnd_output_wire                : std_logic;                     -- Round2resetGND:output -> Round2:reset
	signal multiplexer4user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer4user_aclrGND:output -> Multiplexer4:user_aclr
	signal multiplexer4enavcc_output_wire            : std_logic;                     -- Multiplexer4enaVCC:output -> Multiplexer4:ena
	signal multiplexer1user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire            : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal multiplexer2user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer2user_aclrGND:output -> Multiplexer2:user_aclr
	signal multiplexer2enavcc_output_wire            : std_logic;                     -- Multiplexer2enaVCC:output -> Multiplexer2:ena
	signal rounduser_aclrgnd_output_wire             : std_logic;                     -- Rounduser_aclrGND:output -> Round:user_aclr
	signal roundenavcc_output_wire                   : std_logic;                     -- RoundenaVCC:output -> Round:ena
	signal roundresetgnd_output_wire                 : std_logic;                     -- RoundresetGND:output -> Round:reset
	signal pipelined_adder15user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder15user_aclrGND:output -> Pipelined_Adder15:user_aclr
	signal pipelined_adder15enavcc_output_wire       : std_logic;                     -- Pipelined_Adder15enaVCC:output -> Pipelined_Adder15:ena
	signal pipelined_adder14user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder14user_aclrGND:output -> Pipelined_Adder14:user_aclr
	signal pipelined_adder14enavcc_output_wire       : std_logic;                     -- Pipelined_Adder14enaVCC:output -> Pipelined_Adder14:ena
	signal pipelined_adder13user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder13user_aclrGND:output -> Pipelined_Adder13:user_aclr
	signal pipelined_adder13enavcc_output_wire       : std_logic;                     -- Pipelined_Adder13enaVCC:output -> Pipelined_Adder13:ena
	signal pipelined_adder12user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder12user_aclrGND:output -> Pipelined_Adder12:user_aclr
	signal pipelined_adder12enavcc_output_wire       : std_logic;                     -- Pipelined_Adder12enaVCC:output -> Pipelined_Adder12:ena
	signal pipelined_adder11user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder11user_aclrGND:output -> Pipelined_Adder11:user_aclr
	signal pipelined_adder11enavcc_output_wire       : std_logic;                     -- Pipelined_Adder11enaVCC:output -> Pipelined_Adder11:ena
	signal pipelined_adder10user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder10user_aclrGND:output -> Pipelined_Adder10:user_aclr
	signal pipelined_adder10enavcc_output_wire       : std_logic;                     -- Pipelined_Adder10enaVCC:output -> Pipelined_Adder10:ena
	signal multiplexer7user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer7user_aclrGND:output -> Multiplexer7:user_aclr
	signal multiplexer7enavcc_output_wire            : std_logic;                     -- Multiplexer7enaVCC:output -> Multiplexer7:ena
	signal multiplexer8user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer8user_aclrGND:output -> Multiplexer8:user_aclr
	signal multiplexer8enavcc_output_wire            : std_logic;                     -- Multiplexer8enaVCC:output -> Multiplexer8:ena
	signal multiplexer5user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer5user_aclrGND:output -> Multiplexer5:user_aclr
	signal multiplexer5enavcc_output_wire            : std_logic;                     -- Multiplexer5enaVCC:output -> Multiplexer5:ena
	signal multiplexer6user_aclrgnd_output_wire      : std_logic;                     -- Multiplexer6user_aclrGND:output -> Multiplexer6:user_aclr
	signal multiplexer6enavcc_output_wire            : std_logic;                     -- Multiplexer6enaVCC:output -> Multiplexer6:ena
	signal bus_conversion5_output_wire               : std_logic_vector(12 downto 0); -- Bus_Conversion5:output -> [Comparator1:dataa, Comparator2:datab, Comparator:dataa, Multiplexer1:in0, Multiplexer:in0]
	signal bus_conversion10_output_wire              : std_logic_vector(12 downto 0); -- Bus_Conversion10:output -> [Comparator3:dataa, Comparator4:dataa, Comparator5:datab, Multiplexer3:in0, Multiplexer4:in0]
	signal bus_conversion18_output_wire              : std_logic_vector(12 downto 0); -- Bus_Conversion18:output -> [Comparator6:dataa, Comparator7:dataa, Comparator8:datab, Multiplexer6:in0, Multiplexer7:in0]
	signal multiplexer1_result_wire                  : std_logic_vector(12 downto 0); -- Multiplexer1:result -> Multiplexer2:in0
	signal multiplexer_result_wire                   : std_logic_vector(12 downto 0); -- Multiplexer:result -> Multiplexer2:in1
	signal multiplexer4_result_wire                  : std_logic_vector(12 downto 0); -- Multiplexer4:result -> Multiplexer5:in0
	signal multiplexer3_result_wire                  : std_logic_vector(12 downto 0); -- Multiplexer3:result -> Multiplexer5:in1
	signal multiplexer7_result_wire                  : std_logic_vector(12 downto 0); -- Multiplexer7:result -> Multiplexer8:in0
	signal multiplexer6_result_wire                  : std_logic_vector(12 downto 0); -- Multiplexer6:result -> Multiplexer8:in1
	signal bus_conversion3_output_wire               : std_logic_vector(30 downto 0); -- Bus_Conversion3:output -> Pipelined_Adder1:dataa
	signal bus_conversion1_output_wire               : std_logic_vector(30 downto 0); -- Bus_Conversion1:output -> Pipelined_Adder1:datab
	signal multiplexer5_result_wire                  : std_logic_vector(12 downto 0); -- Multiplexer5:result -> Pipelined_Adder10:dataa
	signal bus_conversion17_output_wire              : std_logic_vector(30 downto 0); -- Bus_Conversion17:output -> Pipelined_Adder11:dataa
	signal bus_conversion11_output_wire              : std_logic_vector(30 downto 0); -- Bus_Conversion11:output -> Pipelined_Adder11:datab
	signal pipelined_adder11_result_wire             : std_logic_vector(30 downto 0); -- Pipelined_Adder11:result -> Pipelined_Adder12:dataa
	signal bus_conversion16_output_wire              : std_logic_vector(30 downto 0); -- Bus_Conversion16:output -> Pipelined_Adder12:datab
	signal pipelined_adder12_result_wire             : std_logic_vector(30 downto 0); -- Pipelined_Adder12:result -> Pipelined_Adder13:dataa
	signal bus_conversion12_output_wire              : std_logic_vector(30 downto 0); -- Bus_Conversion12:output -> Pipelined_Adder13:datab
	signal pipelined_adder13_result_wire             : std_logic_vector(30 downto 0); -- Pipelined_Adder13:result -> Pipelined_Adder14:dataa
	signal bus_conversion15_output_wire              : std_logic_vector(30 downto 0); -- Bus_Conversion15:output -> Pipelined_Adder14:datab
	signal multiplexer8_result_wire                  : std_logic_vector(12 downto 0); -- Multiplexer8:result -> Pipelined_Adder15:dataa
	signal pipelined_adder1_result_wire              : std_logic_vector(30 downto 0); -- Pipelined_Adder1:result -> Pipelined_Adder2:dataa
	signal bus_conversion2_output_wire               : std_logic_vector(30 downto 0); -- Bus_Conversion2:output -> Pipelined_Adder2:datab
	signal bus_conversion9_output_wire               : std_logic_vector(30 downto 0); -- Bus_Conversion9:output -> Pipelined_Adder3:dataa
	signal bus_conversion4_output_wire               : std_logic_vector(30 downto 0); -- Bus_Conversion4:output -> Pipelined_Adder3:datab
	signal pipelined_adder3_result_wire              : std_logic_vector(30 downto 0); -- Pipelined_Adder3:result -> Pipelined_Adder4:dataa
	signal bus_conversion8_output_wire               : std_logic_vector(30 downto 0); -- Bus_Conversion8:output -> Pipelined_Adder4:datab
	signal pipelined_adder4_result_wire              : std_logic_vector(30 downto 0); -- Pipelined_Adder4:result -> Pipelined_Adder5:dataa
	signal bus_conversion6_output_wire               : std_logic_vector(30 downto 0); -- Bus_Conversion6:output -> Pipelined_Adder5:datab
	signal pipelined_adder5_result_wire              : std_logic_vector(30 downto 0); -- Pipelined_Adder5:result -> Pipelined_Adder6:dataa
	signal bus_conversion7_output_wire               : std_logic_vector(30 downto 0); -- Bus_Conversion7:output -> Pipelined_Adder6:datab
	signal pipelined_adder2_result_wire              : std_logic_vector(30 downto 0); -- Pipelined_Adder2:result -> Pipelined_Adder7:dataa
	signal bus_conversion13_output_wire              : std_logic_vector(30 downto 0); -- Bus_Conversion13:output -> Pipelined_Adder7:datab
	signal pipelined_adder7_result_wire              : std_logic_vector(30 downto 0); -- Pipelined_Adder7:result -> Pipelined_Adder8:dataa
	signal bus_conversion14_output_wire              : std_logic_vector(30 downto 0); -- Bus_Conversion14:output -> Pipelined_Adder8:datab
	signal multiplexer2_result_wire                  : std_logic_vector(12 downto 0); -- Multiplexer2:result -> Pipelined_Adder9:dataa
	signal pipelined_adder8_result_wire              : std_logic_vector(30 downto 0); -- Pipelined_Adder8:result -> Round:datain
	signal pipelined_adder6_result_wire              : std_logic_vector(30 downto 0); -- Pipelined_Adder6:result -> Round1:datain
	signal pipelined_adder14_result_wire             : std_logic_vector(30 downto 0); -- Pipelined_Adder14:result -> Round2:datain
	signal un1_output_wire                           : std_logic_vector(12 downto 0); -- Un1:output -> [Comparator:datab, Multiplexer:in1]
	signal un10_output_wire                          : std_logic_vector(12 downto 0); -- Un10:output -> Pipelined_Adder9:datab
	signal un11_output_wire                          : std_logic_vector(12 downto 0); -- Un11:output -> [Comparator7:datab, Multiplexer7:in1]
	signal un2_output_wire                           : std_logic_vector(12 downto 0); -- Un2:output -> [Comparator1:datab, Multiplexer1:in1]
	signal un4_output_wire                           : std_logic_vector(12 downto 0); -- Un4:output -> [Comparator3:datab, Multiplexer3:in1]
	signal un5_output_wire                           : std_logic_vector(12 downto 0); -- Un5:output -> Pipelined_Adder10:datab
	signal un6_output_wire                           : std_logic_vector(12 downto 0); -- Un6:output -> [Comparator4:datab, Multiplexer4:in1]
	signal un8_output_wire                           : std_logic_vector(12 downto 0); -- Un8:output -> [Comparator6:datab, Multiplexer6:in1]
	signal un9_output_wire                           : std_logic_vector(12 downto 0); -- Un9:output -> Pipelined_Adder15:datab
	signal pipelined_adder9_result_wire              : std_logic_vector(12 downto 0); -- Pipelined_Adder9:result -> Vacont_int_0:input
	signal pipelined_adder10_result_wire             : std_logic_vector(12 downto 0); -- Pipelined_Adder10:result -> Vbcont_int_0:input
	signal pipelined_adder15_result_wire             : std_logic_vector(12 downto 0); -- Pipelined_Adder15:result -> Vccont_int_0:input
	signal vbcont_0_output_wire                      : std_logic_vector(13 downto 0); -- vbcont_0:output -> [cast33:input, cast41:input, cast42:input, cast43:input, cast44:input]
	signal cast33_output_wire                        : std_logic_vector(23 downto 0); -- cast33:output -> BinaryPointCasting_x1:input
	signal vccont_0_output_wire                      : std_logic_vector(13 downto 0); -- vccont_0:output -> [cast34:input, cast36:input, cast45:input, cast46:input, cast47:input]
	signal cast34_output_wire                        : std_logic_vector(23 downto 0); -- cast34:output -> BinaryPointCasting_x10:input
	signal vacont_0_output_wire                      : std_logic_vector(13 downto 0); -- vacont_0:output -> [cast35:input, cast37:input, cast38:input, cast39:input, cast40:input]
	signal cast35_output_wire                        : std_logic_vector(23 downto 0); -- cast35:output -> BinaryPointCasting_x1024:input
	signal cast36_output_wire                        : std_logic_vector(23 downto 0); -- cast36:output -> BinaryPointCasting_x11:input
	signal cast37_output_wire                        : std_logic_vector(23 downto 0); -- cast37:output -> BinaryPointCasting_x128:input
	signal cast38_output_wire                        : std_logic_vector(23 downto 0); -- cast38:output -> BinaryPointCasting_x16:input
	signal cast39_output_wire                        : std_logic_vector(23 downto 0); -- cast39:output -> BinaryPointCasting_x2:input
	signal cast40_output_wire                        : std_logic_vector(23 downto 0); -- cast40:output -> BinaryPointCasting_x256:input
	signal cast41_output_wire                        : std_logic_vector(23 downto 0); -- cast41:output -> BinaryPointCasting_x3:input
	signal cast42_output_wire                        : std_logic_vector(23 downto 0); -- cast42:output -> BinaryPointCasting_x4:input
	signal cast43_output_wire                        : std_logic_vector(23 downto 0); -- cast43:output -> BinaryPointCasting_x5:input
	signal cast44_output_wire                        : std_logic_vector(23 downto 0); -- cast44:output -> BinaryPointCasting_x6:input
	signal cast45_output_wire                        : std_logic_vector(23 downto 0); -- cast45:output -> BinaryPointCasting_x7:input
	signal cast46_output_wire                        : std_logic_vector(23 downto 0); -- cast46:output -> BinaryPointCasting_x8:input
	signal cast47_output_wire                        : std_logic_vector(23 downto 0); -- cast47:output -> BinaryPointCasting_x9:input
	signal binarypointcasting_x256_output_wire       : std_logic_vector(23 downto 0); -- BinaryPointCasting_x256:output -> cast48:input
	signal cast48_output_wire                        : std_logic_vector(30 downto 0); -- cast48:output -> Bus_Conversion1:input
	signal binarypointcasting_x11_output_wire        : std_logic_vector(23 downto 0); -- BinaryPointCasting_x11:output -> cast49:input
	signal cast49_output_wire                        : std_logic_vector(30 downto 0); -- cast49:output -> Bus_Conversion11:input
	signal binarypointcasting_x9_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x9:output -> cast50:input
	signal cast50_output_wire                        : std_logic_vector(30 downto 0); -- cast50:output -> Bus_Conversion12:input
	signal binarypointcasting_x16_output_wire        : std_logic_vector(23 downto 0); -- BinaryPointCasting_x16:output -> cast51:input
	signal cast51_output_wire                        : std_logic_vector(30 downto 0); -- cast51:output -> Bus_Conversion13:input
	signal binarypointcasting_x2_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x2:output -> cast52:input
	signal cast52_output_wire                        : std_logic_vector(30 downto 0); -- cast52:output -> Bus_Conversion14:input
	signal binarypointcasting_x10_output_wire        : std_logic_vector(23 downto 0); -- BinaryPointCasting_x10:output -> cast53:input
	signal cast53_output_wire                        : std_logic_vector(30 downto 0); -- cast53:output -> Bus_Conversion15:input
	signal binarypointcasting_x8_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x8:output -> cast54:input
	signal cast54_output_wire                        : std_logic_vector(30 downto 0); -- cast54:output -> Bus_Conversion16:input
	signal binarypointcasting_x7_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x7:output -> cast55:input
	signal cast55_output_wire                        : std_logic_vector(30 downto 0); -- cast55:output -> Bus_Conversion17:input
	signal binarypointcasting_x128_output_wire       : std_logic_vector(23 downto 0); -- BinaryPointCasting_x128:output -> cast56:input
	signal cast56_output_wire                        : std_logic_vector(30 downto 0); -- cast56:output -> Bus_Conversion2:input
	signal binarypointcasting_x1024_output_wire      : std_logic_vector(23 downto 0); -- BinaryPointCasting_x1024:output -> cast57:input
	signal cast57_output_wire                        : std_logic_vector(30 downto 0); -- cast57:output -> Bus_Conversion3:input
	signal binarypointcasting_x6_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x6:output -> cast58:input
	signal cast58_output_wire                        : std_logic_vector(30 downto 0); -- cast58:output -> Bus_Conversion4:input
	signal binarypointcasting_x4_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x4:output -> cast59:input
	signal cast59_output_wire                        : std_logic_vector(30 downto 0); -- cast59:output -> Bus_Conversion6:input
	signal binarypointcasting_x5_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x5:output -> cast60:input
	signal cast60_output_wire                        : std_logic_vector(30 downto 0); -- cast60:output -> Bus_Conversion7:input
	signal binarypointcasting_x3_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x3:output -> cast61:input
	signal cast61_output_wire                        : std_logic_vector(30 downto 0); -- cast61:output -> Bus_Conversion8:input
	signal binarypointcasting_x1_output_wire         : std_logic_vector(23 downto 0); -- BinaryPointCasting_x1:output -> cast62:input
	signal cast62_output_wire                        : std_logic_vector(30 downto 0); -- cast62:output -> Bus_Conversion9:input
	signal comparator_result_wire                    : std_logic;                     -- Comparator:result -> cast63:input
	signal cast63_output_wire                        : std_logic_vector(0 downto 0);  -- cast63:output -> Multiplexer:sel
	signal comparator1_result_wire                   : std_logic;                     -- Comparator1:result -> cast64:input
	signal cast64_output_wire                        : std_logic_vector(0 downto 0);  -- cast64:output -> Multiplexer1:sel
	signal comparator2_result_wire                   : std_logic;                     -- Comparator2:result -> cast65:input
	signal cast65_output_wire                        : std_logic_vector(0 downto 0);  -- cast65:output -> Multiplexer2:sel
	signal comparator3_result_wire                   : std_logic;                     -- Comparator3:result -> cast66:input
	signal cast66_output_wire                        : std_logic_vector(0 downto 0);  -- cast66:output -> Multiplexer3:sel
	signal comparator4_result_wire                   : std_logic;                     -- Comparator4:result -> cast67:input
	signal cast67_output_wire                        : std_logic_vector(0 downto 0);  -- cast67:output -> Multiplexer4:sel
	signal comparator5_result_wire                   : std_logic;                     -- Comparator5:result -> cast68:input
	signal cast68_output_wire                        : std_logic_vector(0 downto 0);  -- cast68:output -> Multiplexer5:sel
	signal comparator6_result_wire                   : std_logic;                     -- Comparator6:result -> cast69:input
	signal cast69_output_wire                        : std_logic_vector(0 downto 0);  -- cast69:output -> Multiplexer6:sel
	signal comparator7_result_wire                   : std_logic;                     -- Comparator7:result -> cast70:input
	signal cast70_output_wire                        : std_logic_vector(0 downto 0);  -- cast70:output -> Multiplexer7:sel
	signal comparator8_result_wire                   : std_logic;                     -- Comparator8:result -> cast71:input
	signal cast71_output_wire                        : std_logic_vector(0 downto 0);  -- cast71:output -> Multiplexer8:sel
	signal round_dataout_wire                        : std_logic_vector(12 downto 0); -- Round:dataout -> cast72:input
	signal cast72_output_wire                        : std_logic_vector(12 downto 0); -- cast72:output -> Bus_Conversion5:input
	signal round1_dataout_wire                       : std_logic_vector(12 downto 0); -- Round1:dataout -> cast73:input
	signal cast73_output_wire                        : std_logic_vector(12 downto 0); -- cast73:output -> Bus_Conversion10:input
	signal round2_dataout_wire                       : std_logic_vector(12 downto 0); -- Round2:dataout -> cast74:input
	signal cast74_output_wire                        : std_logic_vector(12 downto 0); -- cast74:output -> Bus_Conversion18:input
	signal un12_output_wire                          : std_logic_vector(10 downto 0); -- Un12:output -> cast75:input
	signal cast75_output_wire                        : std_logic_vector(12 downto 0); -- cast75:output -> Comparator8:dataa
	signal un3_output_wire                           : std_logic_vector(10 downto 0); -- Un3:output -> cast76:input
	signal cast76_output_wire                        : std_logic_vector(12 downto 0); -- cast76:output -> Comparator2:dataa
	signal un7_output_wire                           : std_logic_vector(10 downto 0); -- Un7:output -> cast77:input
	signal cast77_output_wire                        : std_logic_vector(12 downto 0); -- cast77:output -> Comparator5:dataa
	signal clock_0_clock_output_clk                  : std_logic;                     -- Clock_0:clock_out -> [Comparator1:clock, Comparator2:clock, Comparator3:clock, Comparator4:clock, Comparator5:clock, Comparator6:clock, Comparator7:clock, Comparator8:clock, Comparator:clock, Multiplexer1:clock, Multiplexer2:clock, Multiplexer3:clock, Multiplexer4:clock, Multiplexer5:clock, Multiplexer6:clock, Multiplexer7:clock, Multiplexer8:clock, Multiplexer:clock, Pipelined_Adder10:clock, Pipelined_Adder11:clock, Pipelined_Adder12:clock, Pipelined_Adder13:clock, Pipelined_Adder14:clock, Pipelined_Adder15:clock, Pipelined_Adder1:clock, Pipelined_Adder2:clock, Pipelined_Adder3:clock, Pipelined_Adder4:clock, Pipelined_Adder5:clock, Pipelined_Adder6:clock, Pipelined_Adder7:clock, Pipelined_Adder8:clock, Pipelined_Adder9:clock, Round1:clk, Round2:clk, Round:clk]
	signal clock_0_clock_output_reset                : std_logic;                     -- Clock_0:aclr_out -> [Comparator1:sclr, Comparator2:sclr, Comparator3:sclr, Comparator4:sclr, Comparator5:sclr, Comparator6:sclr, Comparator7:sclr, Comparator8:sclr, Comparator:sclr, Multiplexer1:aclr, Multiplexer2:aclr, Multiplexer3:aclr, Multiplexer4:aclr, Multiplexer5:aclr, Multiplexer6:aclr, Multiplexer7:aclr, Multiplexer8:aclr, Multiplexer:aclr, Pipelined_Adder10:aclr, Pipelined_Adder11:aclr, Pipelined_Adder12:aclr, Pipelined_Adder13:aclr, Pipelined_Adder14:aclr, Pipelined_Adder15:aclr, Pipelined_Adder1:aclr, Pipelined_Adder2:aclr, Pipelined_Adder3:aclr, Pipelined_Adder4:aclr, Pipelined_Adder5:aclr, Pipelined_Adder6:aclr, Pipelined_Adder7:aclr, Pipelined_Adder8:aclr, Pipelined_Adder9:aclr, Round1:reset, Round2:reset, Round:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => cast63_output_wire,                  --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => bus_conversion5_output_wire,         --        in0.wire
			in1       => un1_output_wire                      --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	comparator : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altaleb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,    -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,  --           .reset
			dataa  => bus_conversion5_output_wire, --      dataa.wire
			datab  => un1_output_wire,             --      datab.wire
			result => comparator_result_wire       --     result.wire
		);

	binarypointcasting_x1024 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast35_output_wire,                   --  input.wire
			output => binarypointcasting_x1024_output_wire  -- output.wire
		);

	pipelined_adder9 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 13
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => multiplexer2_result_wire,                 --      dataa.wire
			datab     => un10_output_wire,                         --      datab.wire
			result    => pipelined_adder9_result_wire,             --     result.wire
			user_aclr => pipelined_adder9user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder9enavcc_output_wire        --        ena.wire
		);

	pipelined_adder9user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder9user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder9enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder9enavcc_output_wire  -- output.wire
		);

	pipelined_adder4 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => pipelined_adder3_result_wire,             --      dataa.wire
			datab     => bus_conversion8_output_wire,              --      datab.wire
			result    => pipelined_adder4_result_wire,             --     result.wire
			user_aclr => pipelined_adder4user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder4enavcc_output_wire        --        ena.wire
		);

	pipelined_adder4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder4user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder4enavcc_output_wire  -- output.wire
		);

	un2 : component alt_dspbuilder_constant_GN2SAWFEVT
		generic map (
			BitPattern => "0010110010010",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un2_output_wire  -- output.wire
		);

	pipelined_adder3 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => bus_conversion9_output_wire,              --      dataa.wire
			datab     => bus_conversion4_output_wire,              --      datab.wire
			result    => pipelined_adder3_result_wire,             --     result.wire
			user_aclr => pipelined_adder3user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder3enavcc_output_wire        --        ena.wire
		);

	pipelined_adder3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder3user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder3enavcc_output_wire  -- output.wire
		);

	un1 : component alt_dspbuilder_constant_GNC5QUYE2B
		generic map (
			BitPattern => "1101001101110",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un1_output_wire  -- output.wire
		);

	pipelined_adder2 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => pipelined_adder1_result_wire,             --      dataa.wire
			datab     => bus_conversion2_output_wire,              --      datab.wire
			result    => pipelined_adder2_result_wire,             --     result.wire
			user_aclr => pipelined_adder2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder2enavcc_output_wire        --        ena.wire
		);

	pipelined_adder2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder2user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder2enavcc_output_wire  -- output.wire
		);

	un4 : component alt_dspbuilder_constant_GNC5QUYE2B
		generic map (
			BitPattern => "1101001101110",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un4_output_wire  -- output.wire
		);

	bus_conversion9 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast62_output_wire,          --  input.wire
			output => bus_conversion9_output_wire  -- output.wire
		);

	pipelined_adder1 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => bus_conversion3_output_wire,              --      dataa.wire
			datab     => bus_conversion1_output_wire,              --      datab.wire
			result    => pipelined_adder1_result_wire,             --     result.wire
			user_aclr => pipelined_adder1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder1enavcc_output_wire        --        ena.wire
		);

	pipelined_adder1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder1user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder1enavcc_output_wire  -- output.wire
		);

	un3 : component alt_dspbuilder_constant_GNCOTI3HOF
		generic map (
			BitPattern => "00000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 11
		)
		port map (
			output => un3_output_wire  -- output.wire
		);

	bus_conversion8 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast61_output_wire,          --  input.wire
			output => bus_conversion8_output_wire  -- output.wire
		);

	pipelined_adder8 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => pipelined_adder7_result_wire,             --      dataa.wire
			datab     => bus_conversion14_output_wire,             --      datab.wire
			result    => pipelined_adder8_result_wire,             --     result.wire
			user_aclr => pipelined_adder8user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder8enavcc_output_wire        --        ena.wire
		);

	pipelined_adder8user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder8user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder8enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder8enavcc_output_wire  -- output.wire
		);

	un6 : component alt_dspbuilder_constant_GN2SAWFEVT
		generic map (
			BitPattern => "0010110010010",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un6_output_wire  -- output.wire
		);

	bus_conversion7 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast60_output_wire,          --  input.wire
			output => bus_conversion7_output_wire  -- output.wire
		);

	pipelined_adder7 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => pipelined_adder2_result_wire,             --      dataa.wire
			datab     => bus_conversion13_output_wire,             --      datab.wire
			result    => pipelined_adder7_result_wire,             --     result.wire
			user_aclr => pipelined_adder7user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder7enavcc_output_wire        --        ena.wire
		);

	pipelined_adder7user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder7user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder7enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder7enavcc_output_wire  -- output.wire
		);

	un5 : component alt_dspbuilder_constant_GNGPCXCFCV
		generic map (
			BitPattern => "0011101011111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un5_output_wire  -- output.wire
		);

	bus_conversion6 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast59_output_wire,          --  input.wire
			output => bus_conversion6_output_wire  -- output.wire
		);

	pipelined_adder6 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => pipelined_adder5_result_wire,             --      dataa.wire
			datab     => bus_conversion7_output_wire,              --      datab.wire
			result    => pipelined_adder6_result_wire,             --     result.wire
			user_aclr => pipelined_adder6user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder6enavcc_output_wire        --        ena.wire
		);

	pipelined_adder6user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder6user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder6enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder6enavcc_output_wire  -- output.wire
		);

	un8 : component alt_dspbuilder_constant_GNC5QUYE2B
		generic map (
			BitPattern => "1101001101110",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un8_output_wire  -- output.wire
		);

	bus_conversion5 : component alt_dspbuilder_cast_GNA5AA6QPF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast72_output_wire,          --  input.wire
			output => bus_conversion5_output_wire  -- output.wire
		);

	pipelined_adder5 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => pipelined_adder4_result_wire,             --      dataa.wire
			datab     => bus_conversion6_output_wire,              --      datab.wire
			result    => pipelined_adder5_result_wire,             --     result.wire
			user_aclr => pipelined_adder5user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder5enavcc_output_wire        --        ena.wire
		);

	pipelined_adder5user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder5user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder5enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder5enavcc_output_wire  -- output.wire
		);

	un7 : component alt_dspbuilder_constant_GNCOTI3HOF
		generic map (
			BitPattern => "00000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 11
		)
		port map (
			output => un7_output_wire  -- output.wire
		);

	bus_conversion17 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast55_output_wire,           --  input.wire
			output => bus_conversion17_output_wire  -- output.wire
		);

	bus_conversion4 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast58_output_wire,          --  input.wire
			output => bus_conversion4_output_wire  -- output.wire
		);

	bus_conversion16 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast54_output_wire,           --  input.wire
			output => bus_conversion16_output_wire  -- output.wire
		);

	bus_conversion3 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast57_output_wire,          --  input.wire
			output => bus_conversion3_output_wire  -- output.wire
		);

	un9 : component alt_dspbuilder_constant_GNGPCXCFCV
		generic map (
			BitPattern => "0011101011111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un9_output_wire  -- output.wire
		);

	vccont_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => vccont,               --  input.wire
			output => vccont_0_output_wire  -- output.wire
		);

	bus_conversion15 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast53_output_wire,           --  input.wire
			output => bus_conversion15_output_wire  -- output.wire
		);

	bus_conversion2 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast56_output_wire,          --  input.wire
			output => bus_conversion2_output_wire  -- output.wire
		);

	bus_conversion1 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast48_output_wire,          --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	bus_conversion14 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast52_output_wire,           --  input.wire
			output => bus_conversion14_output_wire  -- output.wire
		);

	vbcont_int_0 : component alt_dspbuilder_port_GNKZFR37ZH
		port map (
			input  => pipelined_adder10_result_wire, --  input.wire
			output => Vbcont_int                     -- output.wire
		);

	bus_conversion18 : component alt_dspbuilder_cast_GNA5AA6QPF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast74_output_wire,           --  input.wire
			output => bus_conversion18_output_wire  -- output.wire
		);

	comparator8 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altageb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,     -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,   --           .reset
			dataa  => cast75_output_wire,           --      dataa.wire
			datab  => bus_conversion18_output_wire, --      datab.wire
			result => comparator8_result_wire       --     result.wire
		);

	comparator7 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altageb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,     -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,   --           .reset
			dataa  => bus_conversion18_output_wire, --      dataa.wire
			datab  => un11_output_wire,             --      datab.wire
			result => comparator7_result_wire       --     result.wire
		);

	comparator6 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altaleb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,     -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,   --           .reset
			dataa  => bus_conversion18_output_wire, --      dataa.wire
			datab  => un8_output_wire,              --      datab.wire
			result => comparator6_result_wire       --     result.wire
		);

	bus_conversion13 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast51_output_wire,           --  input.wire
			output => bus_conversion13_output_wire  -- output.wire
		);

	bus_conversion12 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast50_output_wire,           --  input.wire
			output => bus_conversion12_output_wire  -- output.wire
		);

	bus_conversion11 : component alt_dspbuilder_cast_GN32Z4PX3B
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast49_output_wire,           --  input.wire
			output => bus_conversion11_output_wire  -- output.wire
		);

	bus_conversion10 : component alt_dspbuilder_cast_GNA5AA6QPF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast73_output_wire,           --  input.wire
			output => bus_conversion10_output_wire  -- output.wire
		);

	un10 : component alt_dspbuilder_constant_GNGPCXCFCV
		generic map (
			BitPattern => "0011101011111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un10_output_wire  -- output.wire
		);

	vbcont_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => vbcont,               --  input.wire
			output => vbcont_0_output_wire  -- output.wire
		);

	un11 : component alt_dspbuilder_constant_GN2SAWFEVT
		generic map (
			BitPattern => "0010110010010",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => un11_output_wire  -- output.wire
		);

	un12 : component alt_dspbuilder_constant_GNCOTI3HOF
		generic map (
			BitPattern => "00000000000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 11
		)
		port map (
			output => un12_output_wire  -- output.wire
		);

	vacont_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => vacont,               --  input.wire
			output => vacont_0_output_wire  -- output.wire
		);

	binarypointcasting_x256 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast40_output_wire,                  --  input.wire
			output => binarypointcasting_x256_output_wire  -- output.wire
		);

	round1 : component alt_dspbuilder_round_GNJN4GDIEL
		generic map (
			OUT_WIDTH_g     => 13,
			IN_WIDTH_g      => 31,
			PIPELINE_g      => 0,
			ROUNDING_TYPE_g => "TRUNCATE_LOW",
			SIGNED_g        => 1
		)
		port map (
			clk       => clock_0_clock_output_clk,       -- clk_reset.clk
			reset     => clock_0_clock_output_reset,     --          .reset
			datain    => pipelined_adder6_result_wire,   --    datain.wire
			dataout   => round1_dataout_wire,            --   dataout.wire
			ena       => round1enavcc_output_wire,       --       ena.wire
			user_aclr => round1user_aclrgnd_output_wire  -- user_aclr.wire
		);

	round1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => round1user_aclrgnd_output_wire  -- output.wire
		);

	round1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => round1enavcc_output_wire  -- output.wire
		);

	round1resetgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => round1resetgnd_output_wire  -- output.wire
		);

	multiplexer3 : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast66_output_wire,                   --        sel.wire
			result    => multiplexer3_result_wire,             --     result.wire
			ena       => multiplexer3enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer3user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => bus_conversion10_output_wire,         --        in0.wire
			in1       => un4_output_wire                       --        in1.wire
		);

	multiplexer3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer3user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer3enavcc_output_wire  -- output.wire
		);

	round2 : component alt_dspbuilder_round_GNJN4GDIEL
		generic map (
			OUT_WIDTH_g     => 13,
			IN_WIDTH_g      => 31,
			PIPELINE_g      => 0,
			ROUNDING_TYPE_g => "TRUNCATE_LOW",
			SIGNED_g        => 1
		)
		port map (
			clk       => clock_0_clock_output_clk,       -- clk_reset.clk
			reset     => clock_0_clock_output_reset,     --          .reset
			datain    => pipelined_adder14_result_wire,  --    datain.wire
			dataout   => round2_dataout_wire,            --   dataout.wire
			ena       => round2enavcc_output_wire,       --       ena.wire
			user_aclr => round2user_aclrgnd_output_wire  -- user_aclr.wire
		);

	round2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => round2user_aclrgnd_output_wire  -- output.wire
		);

	round2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => round2enavcc_output_wire  -- output.wire
		);

	round2resetgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => round2resetgnd_output_wire  -- output.wire
		);

	multiplexer4 : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast67_output_wire,                   --        sel.wire
			result    => multiplexer4_result_wire,             --     result.wire
			ena       => multiplexer4enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer4user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => bus_conversion10_output_wire,         --        in0.wire
			in1       => un6_output_wire                       --        in1.wire
		);

	multiplexer4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer4user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer4enavcc_output_wire  -- output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast64_output_wire,                   --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => bus_conversion5_output_wire,          --        in0.wire
			in1       => un2_output_wire                       --        in1.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	multiplexer2 : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast65_output_wire,                   --        sel.wire
			result    => multiplexer2_result_wire,             --     result.wire
			ena       => multiplexer2enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer2user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => multiplexer1_result_wire,             --        in0.wire
			in1       => multiplexer_result_wire               --        in1.wire
		);

	multiplexer2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer2user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer2enavcc_output_wire  -- output.wire
		);

	binarypointcasting_x16 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast38_output_wire,                 --  input.wire
			output => binarypointcasting_x16_output_wire  -- output.wire
		);

	binarypointcasting_x11 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast36_output_wire,                 --  input.wire
			output => binarypointcasting_x11_output_wire  -- output.wire
		);

	comparator1 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altageb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,    -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,  --           .reset
			dataa  => bus_conversion5_output_wire, --      dataa.wire
			datab  => un2_output_wire,             --      datab.wire
			result => comparator1_result_wire      --     result.wire
		);

	binarypointcasting_x10 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast34_output_wire,                 --  input.wire
			output => binarypointcasting_x10_output_wire  -- output.wire
		);

	binarypointcasting_x9 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast47_output_wire,                --  input.wire
			output => binarypointcasting_x9_output_wire  -- output.wire
		);

	binarypointcasting_x7 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast45_output_wire,                --  input.wire
			output => binarypointcasting_x7_output_wire  -- output.wire
		);

	comparator5 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altageb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,     -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,   --           .reset
			dataa  => cast77_output_wire,           --      dataa.wire
			datab  => bus_conversion10_output_wire, --      datab.wire
			result => comparator5_result_wire       --     result.wire
		);

	binarypointcasting_x8 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast46_output_wire,                --  input.wire
			output => binarypointcasting_x8_output_wire  -- output.wire
		);

	comparator4 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altageb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,     -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,   --           .reset
			dataa  => bus_conversion10_output_wire, --      dataa.wire
			datab  => un6_output_wire,              --      datab.wire
			result => comparator4_result_wire       --     result.wire
		);

	binarypointcasting_x5 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast43_output_wire,                --  input.wire
			output => binarypointcasting_x5_output_wire  -- output.wire
		);

	comparator3 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altaleb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,     -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,   --           .reset
			dataa  => bus_conversion10_output_wire, --      dataa.wire
			datab  => un4_output_wire,              --      datab.wire
			result => comparator3_result_wire       --     result.wire
		);

	binarypointcasting_x6 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast44_output_wire,                --  input.wire
			output => binarypointcasting_x6_output_wire  -- output.wire
		);

	comparator2 : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altageb",
			lpm_width => 13
		)
		port map (
			clock  => clock_0_clock_output_clk,    -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset,  --           .reset
			dataa  => cast76_output_wire,          --      dataa.wire
			datab  => bus_conversion5_output_wire, --      datab.wire
			result => comparator2_result_wire      --     result.wire
		);

	binarypointcasting_x3 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast41_output_wire,                --  input.wire
			output => binarypointcasting_x3_output_wire  -- output.wire
		);

	binarypointcasting_x4 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast42_output_wire,                --  input.wire
			output => binarypointcasting_x4_output_wire  -- output.wire
		);

	round : component alt_dspbuilder_round_GNJN4GDIEL
		generic map (
			OUT_WIDTH_g     => 13,
			IN_WIDTH_g      => 31,
			PIPELINE_g      => 0,
			ROUNDING_TYPE_g => "TRUNCATE_LOW",
			SIGNED_g        => 1
		)
		port map (
			clk       => clock_0_clock_output_clk,      -- clk_reset.clk
			reset     => clock_0_clock_output_reset,    --          .reset
			datain    => pipelined_adder8_result_wire,  --    datain.wire
			dataout   => round_dataout_wire,            --   dataout.wire
			ena       => roundenavcc_output_wire,       --       ena.wire
			user_aclr => rounduser_aclrgnd_output_wire  -- user_aclr.wire
		);

	rounduser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => rounduser_aclrgnd_output_wire  -- output.wire
		);

	roundenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => roundenavcc_output_wire  -- output.wire
		);

	roundresetgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => roundresetgnd_output_wire  -- output.wire
		);

	binarypointcasting_x1 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast33_output_wire,                --  input.wire
			output => binarypointcasting_x1_output_wire  -- output.wire
		);

	binarypointcasting_x2 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast39_output_wire,                --  input.wire
			output => binarypointcasting_x2_output_wire  -- output.wire
		);

	vccont_int_0 : component alt_dspbuilder_port_GNKZFR37ZH
		port map (
			input  => pipelined_adder15_result_wire, --  input.wire
			output => Vccont_int                     -- output.wire
		);

	pipelined_adder15 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 13
		)
		port map (
			clock     => clock_0_clock_output_clk,                  -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                --           .reset
			dataa     => multiplexer8_result_wire,                  --      dataa.wire
			datab     => un9_output_wire,                           --      datab.wire
			result    => pipelined_adder15_result_wire,             --     result.wire
			user_aclr => pipelined_adder15user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder15enavcc_output_wire        --        ena.wire
		);

	pipelined_adder15user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder15user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder15enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder15enavcc_output_wire  -- output.wire
		);

	pipelined_adder14 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                  -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                --           .reset
			dataa     => pipelined_adder13_result_wire,             --      dataa.wire
			datab     => bus_conversion15_output_wire,              --      datab.wire
			result    => pipelined_adder14_result_wire,             --     result.wire
			user_aclr => pipelined_adder14user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder14enavcc_output_wire        --        ena.wire
		);

	pipelined_adder14user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder14user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder14enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder14enavcc_output_wire  -- output.wire
		);

	vacont_int_0 : component alt_dspbuilder_port_GNKZFR37ZH
		port map (
			input  => pipelined_adder9_result_wire, --  input.wire
			output => Vacont_int                    -- output.wire
		);

	pipelined_adder13 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                  -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                --           .reset
			dataa     => pipelined_adder12_result_wire,             --      dataa.wire
			datab     => bus_conversion12_output_wire,              --      datab.wire
			result    => pipelined_adder13_result_wire,             --     result.wire
			user_aclr => pipelined_adder13user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder13enavcc_output_wire        --        ena.wire
		);

	pipelined_adder13user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder13user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder13enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder13enavcc_output_wire  -- output.wire
		);

	pipelined_adder12 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                  -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                --           .reset
			dataa     => pipelined_adder11_result_wire,             --      dataa.wire
			datab     => bus_conversion16_output_wire,              --      datab.wire
			result    => pipelined_adder12_result_wire,             --     result.wire
			user_aclr => pipelined_adder12user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder12enavcc_output_wire        --        ena.wire
		);

	pipelined_adder12user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder12user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder12enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder12enavcc_output_wire  -- output.wire
		);

	pipelined_adder11 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 31
		)
		port map (
			clock     => clock_0_clock_output_clk,                  -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                --           .reset
			dataa     => bus_conversion17_output_wire,              --      dataa.wire
			datab     => bus_conversion11_output_wire,              --      datab.wire
			result    => pipelined_adder11_result_wire,             --     result.wire
			user_aclr => pipelined_adder11user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder11enavcc_output_wire        --        ena.wire
		);

	pipelined_adder11user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder11user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder11enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder11enavcc_output_wire  -- output.wire
		);

	binarypointcasting_x128 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast37_output_wire,                  --  input.wire
			output => binarypointcasting_x128_output_wire  -- output.wire
		);

	pipelined_adder10 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 13
		)
		port map (
			clock     => clock_0_clock_output_clk,                  -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                --           .reset
			dataa     => multiplexer5_result_wire,                  --      dataa.wire
			datab     => un5_output_wire,                           --      datab.wire
			result    => pipelined_adder10_result_wire,             --     result.wire
			user_aclr => pipelined_adder10user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder10enavcc_output_wire        --        ena.wire
		);

	pipelined_adder10user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder10user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder10enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder10enavcc_output_wire  -- output.wire
		);

	multiplexer7 : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast70_output_wire,                   --        sel.wire
			result    => multiplexer7_result_wire,             --     result.wire
			ena       => multiplexer7enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer7user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => bus_conversion18_output_wire,         --        in0.wire
			in1       => un11_output_wire                      --        in1.wire
		);

	multiplexer7user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer7user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer7enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer7enavcc_output_wire  -- output.wire
		);

	multiplexer8 : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast71_output_wire,                   --        sel.wire
			result    => multiplexer8_result_wire,             --     result.wire
			ena       => multiplexer8enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer8user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => multiplexer7_result_wire,             --        in0.wire
			in1       => multiplexer6_result_wire              --        in1.wire
		);

	multiplexer8user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer8user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer8enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer8enavcc_output_wire  -- output.wire
		);

	multiplexer5 : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast68_output_wire,                   --        sel.wire
			result    => multiplexer5_result_wire,             --     result.wire
			ena       => multiplexer5enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer5user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => multiplexer4_result_wire,             --        in0.wire
			in1       => multiplexer3_result_wire              --        in1.wire
		);

	multiplexer5user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer5user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer5enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer5enavcc_output_wire  -- output.wire
		);

	multiplexer6 : component alt_dspbuilder_multiplexer_GNBGHTTLA2
		generic map (
			number_inputs          => 2,
			pipeline               => 1,
			width                  => 13,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast69_output_wire,                   --        sel.wire
			result    => multiplexer6_result_wire,             --     result.wire
			ena       => multiplexer6enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer6user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => bus_conversion18_output_wire,         --        in0.wire
			in1       => un8_output_wire                       --        in1.wire
		);

	multiplexer6user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer6user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer6enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer6enavcc_output_wire  -- output.wire
		);

	cast33 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vbcont_0_output_wire, --  input.wire
			output => cast33_output_wire    -- output.wire
		);

	cast34 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vccont_0_output_wire, --  input.wire
			output => cast34_output_wire    -- output.wire
		);

	cast35 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vacont_0_output_wire, --  input.wire
			output => cast35_output_wire    -- output.wire
		);

	cast36 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vccont_0_output_wire, --  input.wire
			output => cast36_output_wire    -- output.wire
		);

	cast37 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vacont_0_output_wire, --  input.wire
			output => cast37_output_wire    -- output.wire
		);

	cast38 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vacont_0_output_wire, --  input.wire
			output => cast38_output_wire    -- output.wire
		);

	cast39 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vacont_0_output_wire, --  input.wire
			output => cast39_output_wire    -- output.wire
		);

	cast40 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vacont_0_output_wire, --  input.wire
			output => cast40_output_wire    -- output.wire
		);

	cast41 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vbcont_0_output_wire, --  input.wire
			output => cast41_output_wire    -- output.wire
		);

	cast42 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vbcont_0_output_wire, --  input.wire
			output => cast42_output_wire    -- output.wire
		);

	cast43 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vbcont_0_output_wire, --  input.wire
			output => cast43_output_wire    -- output.wire
		);

	cast44 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vbcont_0_output_wire, --  input.wire
			output => cast44_output_wire    -- output.wire
		);

	cast45 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vccont_0_output_wire, --  input.wire
			output => cast45_output_wire    -- output.wire
		);

	cast46 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vccont_0_output_wire, --  input.wire
			output => cast46_output_wire    -- output.wire
		);

	cast47 : component alt_dspbuilder_cast_GNVPCKFRV6
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vccont_0_output_wire, --  input.wire
			output => cast47_output_wire    -- output.wire
		);

	cast48 : component alt_dspbuilder_cast_GNL533AQU2
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x256_output_wire, --  input.wire
			output => cast48_output_wire                   -- output.wire
		);

	cast49 : component alt_dspbuilder_cast_GNL533AQU2
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x11_output_wire, --  input.wire
			output => cast49_output_wire                  -- output.wire
		);

	cast50 : component alt_dspbuilder_cast_GNSQKJ6AEZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x9_output_wire, --  input.wire
			output => cast50_output_wire                 -- output.wire
		);

	cast51 : component alt_dspbuilder_cast_GNSQKJ6AEZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x16_output_wire, --  input.wire
			output => cast51_output_wire                  -- output.wire
		);

	cast52 : component alt_dspbuilder_cast_GND23XTBOL
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x2_output_wire, --  input.wire
			output => cast52_output_wire                 -- output.wire
		);

	cast53 : component alt_dspbuilder_cast_GND23XTBOL
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x10_output_wire, --  input.wire
			output => cast53_output_wire                  -- output.wire
		);

	cast54 : component alt_dspbuilder_cast_GNRYH7CSLF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x8_output_wire, --  input.wire
			output => cast54_output_wire                 -- output.wire
		);

	cast55 : component alt_dspbuilder_cast_GND5VHVYOD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x7_output_wire, --  input.wire
			output => cast55_output_wire                 -- output.wire
		);

	cast56 : component alt_dspbuilder_cast_GNRYH7CSLF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x128_output_wire, --  input.wire
			output => cast56_output_wire                   -- output.wire
		);

	cast57 : component alt_dspbuilder_cast_GND5VHVYOD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x1024_output_wire, --  input.wire
			output => cast57_output_wire                    -- output.wire
		);

	cast58 : component alt_dspbuilder_cast_GNL533AQU2
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x6_output_wire, --  input.wire
			output => cast58_output_wire                 -- output.wire
		);

	cast59 : component alt_dspbuilder_cast_GNSQKJ6AEZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x4_output_wire, --  input.wire
			output => cast59_output_wire                 -- output.wire
		);

	cast60 : component alt_dspbuilder_cast_GND23XTBOL
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x5_output_wire, --  input.wire
			output => cast60_output_wire                 -- output.wire
		);

	cast61 : component alt_dspbuilder_cast_GNRYH7CSLF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x3_output_wire, --  input.wire
			output => cast61_output_wire                 -- output.wire
		);

	cast62 : component alt_dspbuilder_cast_GND5VHVYOD
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binarypointcasting_x1_output_wire, --  input.wire
			output => cast62_output_wire                 -- output.wire
		);

	cast63 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator_result_wire, --  input.wire
			output => cast63_output_wire      -- output.wire
		);

	cast64 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator1_result_wire, --  input.wire
			output => cast64_output_wire       -- output.wire
		);

	cast65 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator2_result_wire, --  input.wire
			output => cast65_output_wire       -- output.wire
		);

	cast66 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator3_result_wire, --  input.wire
			output => cast66_output_wire       -- output.wire
		);

	cast67 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator4_result_wire, --  input.wire
			output => cast67_output_wire       -- output.wire
		);

	cast68 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator5_result_wire, --  input.wire
			output => cast68_output_wire       -- output.wire
		);

	cast69 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator6_result_wire, --  input.wire
			output => cast69_output_wire       -- output.wire
		);

	cast70 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator7_result_wire, --  input.wire
			output => cast70_output_wire       -- output.wire
		);

	cast71 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator8_result_wire, --  input.wire
			output => cast71_output_wire       -- output.wire
		);

	cast72 : component alt_dspbuilder_cast_GNA5AA6QPF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => round_dataout_wire, --  input.wire
			output => cast72_output_wire  -- output.wire
		);

	cast73 : component alt_dspbuilder_cast_GNA5AA6QPF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => round1_dataout_wire, --  input.wire
			output => cast73_output_wire   -- output.wire
		);

	cast74 : component alt_dspbuilder_cast_GNA5AA6QPF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => round2_dataout_wire, --  input.wire
			output => cast74_output_wire   -- output.wire
		);

	cast75 : component alt_dspbuilder_cast_GNWF56JAW3
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => un12_output_wire,   --  input.wire
			output => cast75_output_wire  -- output.wire
		);

	cast76 : component alt_dspbuilder_cast_GNWF56JAW3
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => un3_output_wire,    --  input.wire
			output => cast76_output_wire  -- output.wire
		);

	cast77 : component alt_dspbuilder_cast_GNWF56JAW3
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => un7_output_wire,    --  input.wire
			output => cast77_output_wire  -- output.wire
		);

end architecture rtl; -- of mem_GN_mem_Conversion_Ioxcont_Int
